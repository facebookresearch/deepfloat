// Copyright (c) Facebook, Inc. and its affiliates. All Rights Reserved.
// All rights reserved.
//
// This source code is licensed under the license found in the
// LICENSE file in the root directory of this source tree.

package Comparison;
  typedef enum { EQ, NE, LT, LE, GT, GE } Type;
endpackage
