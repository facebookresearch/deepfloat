// Copyright (c) Facebook, Inc. and its affiliates. All Rights Reserved.
// All rights reserved.
//
// This source code is licensed under the license found in the
// LICENSE file in the root directory of this source tree.


module Log2LUT_9x8
  (input [8:0] in,
   output logic [8:0] out);

  always_comb begin
    case (in)
      9'b000000000: out = 9'b000000000;
      9'b000000001: out = 9'b000000001;
      9'b000000010: out = 9'b000000001; // overlap
      9'b000000011: out = 9'b000000010;
      9'b000000100: out = 9'b000000011;
      9'b000000101: out = 9'b000000100;
      9'b000000110: out = 9'b000000100; // overlap
      9'b000000111: out = 9'b000000101;
      9'b000001000: out = 9'b000000110;
      9'b000001001: out = 9'b000000110; // overlap
      9'b000001010: out = 9'b000000111;
      9'b000001011: out = 9'b000001000;
      9'b000001100: out = 9'b000001001;
      9'b000001101: out = 9'b000001001; // overlap
      9'b000001110: out = 9'b000001010;
      9'b000001111: out = 9'b000001011;
      9'b000010000: out = 9'b000001011; // overlap
      9'b000010001: out = 9'b000001100;
      9'b000010010: out = 9'b000001101;
      9'b000010011: out = 9'b000001101; // overlap
      9'b000010100: out = 9'b000001110;
      9'b000010101: out = 9'b000001111;
      9'b000010110: out = 9'b000010000;
      9'b000010111: out = 9'b000010000; // overlap
      9'b000011000: out = 9'b000010001;
      9'b000011001: out = 9'b000010010;
      9'b000011010: out = 9'b000010010; // overlap
      9'b000011011: out = 9'b000010011;
      9'b000011100: out = 9'b000010100;
      9'b000011101: out = 9'b000010100; // overlap
      9'b000011110: out = 9'b000010101;
      9'b000011111: out = 9'b000010110;
      9'b000100000: out = 9'b000010110; // overlap
      9'b000100001: out = 9'b000010111;
      9'b000100010: out = 9'b000011000;
      9'b000100011: out = 9'b000011000; // overlap
      9'b000100100: out = 9'b000011001;
      9'b000100101: out = 9'b000011010;
      9'b000100110: out = 9'b000011010; // overlap
      9'b000100111: out = 9'b000011011;
      9'b000101000: out = 9'b000011100;
      9'b000101001: out = 9'b000011100; // overlap
      9'b000101010: out = 9'b000011101;
      9'b000101011: out = 9'b000011110;
      9'b000101100: out = 9'b000011110; // overlap
      9'b000101101: out = 9'b000011111;
      9'b000101110: out = 9'b000100000;
      9'b000101111: out = 9'b000100000; // overlap
      9'b000110000: out = 9'b000100001;
      9'b000110001: out = 9'b000100010;
      9'b000110010: out = 9'b000100010; // overlap
      9'b000110011: out = 9'b000100011;
      9'b000110100: out = 9'b000100100;
      9'b000110101: out = 9'b000100100; // overlap
      9'b000110110: out = 9'b000100101;
      9'b000110111: out = 9'b000100110;
      9'b000111000: out = 9'b000100110; // overlap
      9'b000111001: out = 9'b000100111;
      9'b000111010: out = 9'b000101000;
      9'b000111011: out = 9'b000101000; // overlap
      9'b000111100: out = 9'b000101001;
      9'b000111101: out = 9'b000101010;
      9'b000111110: out = 9'b000101010; // overlap
      9'b000111111: out = 9'b000101011;
      9'b001000000: out = 9'b000101100;
      9'b001000001: out = 9'b000101100; // overlap
      9'b001000010: out = 9'b000101101;
      9'b001000011: out = 9'b000101101; // overlap
      9'b001000100: out = 9'b000101110;
      9'b001000101: out = 9'b000101111;
      9'b001000110: out = 9'b000101111; // overlap
      9'b001000111: out = 9'b000110000;
      9'b001001000: out = 9'b000110001;
      9'b001001001: out = 9'b000110001; // overlap
      9'b001001010: out = 9'b000110010;
      9'b001001011: out = 9'b000110010; // overlap
      9'b001001100: out = 9'b000110011;
      9'b001001101: out = 9'b000110100;
      9'b001001110: out = 9'b000110100; // overlap
      9'b001001111: out = 9'b000110101;
      9'b001010000: out = 9'b000110110;
      9'b001010001: out = 9'b000110110; // overlap
      9'b001010010: out = 9'b000110111;
      9'b001010011: out = 9'b000110111; // overlap
      9'b001010100: out = 9'b000111000;
      9'b001010101: out = 9'b000111001;
      9'b001010110: out = 9'b000111001; // overlap
      9'b001010111: out = 9'b000111010;
      9'b001011000: out = 9'b000111011;
      9'b001011001: out = 9'b000111011; // overlap
      9'b001011010: out = 9'b000111100;
      9'b001011011: out = 9'b000111100; // overlap
      9'b001011100: out = 9'b000111101;
      9'b001011101: out = 9'b000111110;
      9'b001011110: out = 9'b000111110; // overlap
      9'b001011111: out = 9'b000111111;
      9'b001100000: out = 9'b000111111; // overlap
      9'b001100001: out = 9'b001000000;
      9'b001100010: out = 9'b001000001;
      9'b001100011: out = 9'b001000001; // overlap
      9'b001100100: out = 9'b001000010;
      9'b001100101: out = 9'b001000010; // overlap
      9'b001100110: out = 9'b001000011;
      9'b001100111: out = 9'b001000100;
      9'b001101000: out = 9'b001000100; // overlap
      9'b001101001: out = 9'b001000101;
      9'b001101010: out = 9'b001000101; // overlap
      9'b001101011: out = 9'b001000110;
      9'b001101100: out = 9'b001000111;
      9'b001101101: out = 9'b001000111; // overlap
      9'b001101110: out = 9'b001001000;
      9'b001101111: out = 9'b001001000; // overlap
      9'b001110000: out = 9'b001001001;
      9'b001110001: out = 9'b001001010;
      9'b001110010: out = 9'b001001010; // overlap
      9'b001110011: out = 9'b001001011;
      9'b001110100: out = 9'b001001011; // overlap
      9'b001110101: out = 9'b001001100;
      9'b001110110: out = 9'b001001101;
      9'b001110111: out = 9'b001001101; // overlap
      9'b001111000: out = 9'b001001110;
      9'b001111001: out = 9'b001001110; // overlap
      9'b001111010: out = 9'b001001111;
      9'b001111011: out = 9'b001010000;
      9'b001111100: out = 9'b001010000; // overlap
      9'b001111101: out = 9'b001010001;
      9'b001111110: out = 9'b001010001; // overlap
      9'b001111111: out = 9'b001010010;
      9'b010000000: out = 9'b001010010; // overlap
      9'b010000001: out = 9'b001010011;
      9'b010000010: out = 9'b001010100;
      9'b010000011: out = 9'b001010100; // overlap
      9'b010000100: out = 9'b001010101;
      9'b010000101: out = 9'b001010101; // overlap
      9'b010000110: out = 9'b001010110;
      9'b010000111: out = 9'b001010110; // overlap
      9'b010001000: out = 9'b001010111;
      9'b010001001: out = 9'b001011000;
      9'b010001010: out = 9'b001011000; // overlap
      9'b010001011: out = 9'b001011001;
      9'b010001100: out = 9'b001011001; // overlap
      9'b010001101: out = 9'b001011010;
      9'b010001110: out = 9'b001011010; // overlap
      9'b010001111: out = 9'b001011011;
      9'b010010000: out = 9'b001011100;
      9'b010010001: out = 9'b001011100; // overlap
      9'b010010010: out = 9'b001011101;
      9'b010010011: out = 9'b001011101; // overlap
      9'b010010100: out = 9'b001011110;
      9'b010010101: out = 9'b001011110; // overlap
      9'b010010110: out = 9'b001011111;
      9'b010010111: out = 9'b001011111; // overlap
      9'b010011000: out = 9'b001100000;
      9'b010011001: out = 9'b001100001;
      9'b010011010: out = 9'b001100001; // overlap
      9'b010011011: out = 9'b001100010;
      9'b010011100: out = 9'b001100010; // overlap
      9'b010011101: out = 9'b001100011;
      9'b010011110: out = 9'b001100011; // overlap
      9'b010011111: out = 9'b001100100;
      9'b010100000: out = 9'b001100100; // overlap
      9'b010100001: out = 9'b001100101;
      9'b010100010: out = 9'b001100110;
      9'b010100011: out = 9'b001100110; // overlap
      9'b010100100: out = 9'b001100111;
      9'b010100101: out = 9'b001100111; // overlap
      9'b010100110: out = 9'b001101000;
      9'b010100111: out = 9'b001101000; // overlap
      9'b010101000: out = 9'b001101001;
      9'b010101001: out = 9'b001101001; // overlap
      9'b010101010: out = 9'b001101010;
      9'b010101011: out = 9'b001101010; // overlap
      9'b010101100: out = 9'b001101011;
      9'b010101101: out = 9'b001101100;
      9'b010101110: out = 9'b001101100; // overlap
      9'b010101111: out = 9'b001101101;
      9'b010110000: out = 9'b001101101; // overlap
      9'b010110001: out = 9'b001101110;
      9'b010110010: out = 9'b001101110; // overlap
      9'b010110011: out = 9'b001101111;
      9'b010110100: out = 9'b001101111; // overlap
      9'b010110101: out = 9'b001110000;
      9'b010110110: out = 9'b001110000; // overlap
      9'b010110111: out = 9'b001110001;
      9'b010111000: out = 9'b001110001; // overlap
      9'b010111001: out = 9'b001110010;
      9'b010111010: out = 9'b001110010; // overlap
      9'b010111011: out = 9'b001110011;
      9'b010111100: out = 9'b001110100;
      9'b010111101: out = 9'b001110100; // overlap
      9'b010111110: out = 9'b001110101;
      9'b010111111: out = 9'b001110101; // overlap
      9'b011000000: out = 9'b001110110;
      9'b011000001: out = 9'b001110110; // overlap
      9'b011000010: out = 9'b001110111;
      9'b011000011: out = 9'b001110111; // overlap
      9'b011000100: out = 9'b001111000;
      9'b011000101: out = 9'b001111000; // overlap
      9'b011000110: out = 9'b001111001;
      9'b011000111: out = 9'b001111001; // overlap
      9'b011001000: out = 9'b001111010;
      9'b011001001: out = 9'b001111010; // overlap
      9'b011001010: out = 9'b001111011;
      9'b011001011: out = 9'b001111011; // overlap
      9'b011001100: out = 9'b001111100;
      9'b011001101: out = 9'b001111100; // overlap
      9'b011001110: out = 9'b001111101;
      9'b011001111: out = 9'b001111101; // overlap
      9'b011010000: out = 9'b001111110;
      9'b011010001: out = 9'b001111110; // overlap
      9'b011010010: out = 9'b001111111;
      9'b011010011: out = 9'b001111111; // overlap
      9'b011010100: out = 9'b010000000;
      9'b011010101: out = 9'b010000000; // overlap
      9'b011010110: out = 9'b010000001;
      9'b011010111: out = 9'b010000001; // overlap
      9'b011011000: out = 9'b010000010;
      9'b011011001: out = 9'b010000011;
      9'b011011010: out = 9'b010000011; // overlap
      9'b011011011: out = 9'b010000100;
      9'b011011100: out = 9'b010000100; // overlap
      9'b011011101: out = 9'b010000101;
      9'b011011110: out = 9'b010000101; // overlap
      9'b011011111: out = 9'b010000110;
      9'b011100000: out = 9'b010000110; // overlap
      9'b011100001: out = 9'b010000111;
      9'b011100010: out = 9'b010000111; // overlap
      9'b011100011: out = 9'b010001000;
      9'b011100100: out = 9'b010001000; // overlap
      9'b011100101: out = 9'b010001001;
      9'b011100110: out = 9'b010001001; // overlap
      9'b011100111: out = 9'b010001010;
      9'b011101000: out = 9'b010001010; // overlap
      9'b011101001: out = 9'b010001011;
      9'b011101010: out = 9'b010001011; // overlap
      9'b011101011: out = 9'b010001100;
      9'b011101100: out = 9'b010001100; // overlap
      9'b011101101: out = 9'b010001100; // overlap
      9'b011101110: out = 9'b010001101;
      9'b011101111: out = 9'b010001101; // overlap
      9'b011110000: out = 9'b010001110;
      9'b011110001: out = 9'b010001110; // overlap
      9'b011110010: out = 9'b010001111;
      9'b011110011: out = 9'b010001111; // overlap
      9'b011110100: out = 9'b010010000;
      9'b011110101: out = 9'b010010000; // overlap
      9'b011110110: out = 9'b010010001;
      9'b011110111: out = 9'b010010001; // overlap
      9'b011111000: out = 9'b010010010;
      9'b011111001: out = 9'b010010010; // overlap
      9'b011111010: out = 9'b010010011;
      9'b011111011: out = 9'b010010011; // overlap
      9'b011111100: out = 9'b010010100;
      9'b011111101: out = 9'b010010100; // overlap
      9'b011111110: out = 9'b010010101;
      9'b011111111: out = 9'b010010101; // overlap
      9'b100000000: out = 9'b010010110;
      9'b100000001: out = 9'b010010110; // overlap
      9'b100000010: out = 9'b010010111;
      9'b100000011: out = 9'b010010111; // overlap
      9'b100000100: out = 9'b010011000;
      9'b100000101: out = 9'b010011000; // overlap
      9'b100000110: out = 9'b010011001;
      9'b100000111: out = 9'b010011001; // overlap
      9'b100001000: out = 9'b010011010;
      9'b100001001: out = 9'b010011010; // overlap
      9'b100001010: out = 9'b010011011;
      9'b100001011: out = 9'b010011011; // overlap
      9'b100001100: out = 9'b010011011; // overlap
      9'b100001101: out = 9'b010011100;
      9'b100001110: out = 9'b010011100; // overlap
      9'b100001111: out = 9'b010011101;
      9'b100010000: out = 9'b010011101; // overlap
      9'b100010001: out = 9'b010011110;
      9'b100010010: out = 9'b010011110; // overlap
      9'b100010011: out = 9'b010011111;
      9'b100010100: out = 9'b010011111; // overlap
      9'b100010101: out = 9'b010100000;
      9'b100010110: out = 9'b010100000; // overlap
      9'b100010111: out = 9'b010100001;
      9'b100011000: out = 9'b010100001; // overlap
      9'b100011001: out = 9'b010100010;
      9'b100011010: out = 9'b010100010; // overlap
      9'b100011011: out = 9'b010100011;
      9'b100011100: out = 9'b010100011; // overlap
      9'b100011101: out = 9'b010100011; // overlap
      9'b100011110: out = 9'b010100100;
      9'b100011111: out = 9'b010100100; // overlap
      9'b100100000: out = 9'b010100101;
      9'b100100001: out = 9'b010100101; // overlap
      9'b100100010: out = 9'b010100110;
      9'b100100011: out = 9'b010100110; // overlap
      9'b100100100: out = 9'b010100111;
      9'b100100101: out = 9'b010100111; // overlap
      9'b100100110: out = 9'b010101000;
      9'b100100111: out = 9'b010101000; // overlap
      9'b100101000: out = 9'b010101001;
      9'b100101001: out = 9'b010101001; // overlap
      9'b100101010: out = 9'b010101001; // overlap
      9'b100101011: out = 9'b010101010;
      9'b100101100: out = 9'b010101010; // overlap
      9'b100101101: out = 9'b010101011;
      9'b100101110: out = 9'b010101011; // overlap
      9'b100101111: out = 9'b010101100;
      9'b100110000: out = 9'b010101100; // overlap
      9'b100110001: out = 9'b010101101;
      9'b100110010: out = 9'b010101101; // overlap
      9'b100110011: out = 9'b010101101; // overlap
      9'b100110100: out = 9'b010101110;
      9'b100110101: out = 9'b010101110; // overlap
      9'b100110110: out = 9'b010101111;
      9'b100110111: out = 9'b010101111; // overlap
      9'b100111000: out = 9'b010110000;
      9'b100111001: out = 9'b010110000; // overlap
      9'b100111010: out = 9'b010110001;
      9'b100111011: out = 9'b010110001; // overlap
      9'b100111100: out = 9'b010110010;
      9'b100111101: out = 9'b010110010; // overlap
      9'b100111110: out = 9'b010110010; // overlap
      9'b100111111: out = 9'b010110011;
      9'b101000000: out = 9'b010110011; // overlap
      9'b101000001: out = 9'b010110100;
      9'b101000010: out = 9'b010110100; // overlap
      9'b101000011: out = 9'b010110101;
      9'b101000100: out = 9'b010110101; // overlap
      9'b101000101: out = 9'b010110110;
      9'b101000110: out = 9'b010110110; // overlap
      9'b101000111: out = 9'b010110110; // overlap
      9'b101001000: out = 9'b010110111;
      9'b101001001: out = 9'b010110111; // overlap
      9'b101001010: out = 9'b010111000;
      9'b101001011: out = 9'b010111000; // overlap
      9'b101001100: out = 9'b010111001;
      9'b101001101: out = 9'b010111001; // overlap
      9'b101001110: out = 9'b010111001; // overlap
      9'b101001111: out = 9'b010111010;
      9'b101010000: out = 9'b010111010; // overlap
      9'b101010001: out = 9'b010111011;
      9'b101010010: out = 9'b010111011; // overlap
      9'b101010011: out = 9'b010111100;
      9'b101010100: out = 9'b010111100; // overlap
      9'b101010101: out = 9'b010111101;
      9'b101010110: out = 9'b010111101; // overlap
      9'b101010111: out = 9'b010111101; // overlap
      9'b101011000: out = 9'b010111110;
      9'b101011001: out = 9'b010111110; // overlap
      9'b101011010: out = 9'b010111111;
      9'b101011011: out = 9'b010111111; // overlap
      9'b101011100: out = 9'b011000000;
      9'b101011101: out = 9'b011000000; // overlap
      9'b101011110: out = 9'b011000000; // overlap
      9'b101011111: out = 9'b011000001;
      9'b101100000: out = 9'b011000001; // overlap
      9'b101100001: out = 9'b011000010;
      9'b101100010: out = 9'b011000010; // overlap
      9'b101100011: out = 9'b011000011;
      9'b101100100: out = 9'b011000011; // overlap
      9'b101100101: out = 9'b011000011; // overlap
      9'b101100110: out = 9'b011000100;
      9'b101100111: out = 9'b011000100; // overlap
      9'b101101000: out = 9'b011000101;
      9'b101101001: out = 9'b011000101; // overlap
      9'b101101010: out = 9'b011000110;
      9'b101101011: out = 9'b011000110; // overlap
      9'b101101100: out = 9'b011000110; // overlap
      9'b101101101: out = 9'b011000111;
      9'b101101110: out = 9'b011000111; // overlap
      9'b101101111: out = 9'b011001000;
      9'b101110000: out = 9'b011001000; // overlap
      9'b101110001: out = 9'b011001000; // overlap
      9'b101110010: out = 9'b011001001;
      9'b101110011: out = 9'b011001001; // overlap
      9'b101110100: out = 9'b011001010;
      9'b101110101: out = 9'b011001010; // overlap
      9'b101110110: out = 9'b011001011;
      9'b101110111: out = 9'b011001011; // overlap
      9'b101111000: out = 9'b011001011; // overlap
      9'b101111001: out = 9'b011001100;
      9'b101111010: out = 9'b011001100; // overlap
      9'b101111011: out = 9'b011001101;
      9'b101111100: out = 9'b011001101; // overlap
      9'b101111101: out = 9'b011001101; // overlap
      9'b101111110: out = 9'b011001110;
      9'b101111111: out = 9'b011001110; // overlap
      9'b110000000: out = 9'b011001111;
      9'b110000001: out = 9'b011001111; // overlap
      9'b110000010: out = 9'b011010000;
      9'b110000011: out = 9'b011010000; // overlap
      9'b110000100: out = 9'b011010000; // overlap
      9'b110000101: out = 9'b011010001;
      9'b110000110: out = 9'b011010001; // overlap
      9'b110000111: out = 9'b011010010;
      9'b110001000: out = 9'b011010010; // overlap
      9'b110001001: out = 9'b011010010; // overlap
      9'b110001010: out = 9'b011010011;
      9'b110001011: out = 9'b011010011; // overlap
      9'b110001100: out = 9'b011010100;
      9'b110001101: out = 9'b011010100; // overlap
      9'b110001110: out = 9'b011010100; // overlap
      9'b110001111: out = 9'b011010101;
      9'b110010000: out = 9'b011010101; // overlap
      9'b110010001: out = 9'b011010110;
      9'b110010010: out = 9'b011010110; // overlap
      9'b110010011: out = 9'b011010110; // overlap
      9'b110010100: out = 9'b011010111;
      9'b110010101: out = 9'b011010111; // overlap
      9'b110010110: out = 9'b011011000;
      9'b110010111: out = 9'b011011000; // overlap
      9'b110011000: out = 9'b011011000; // overlap
      9'b110011001: out = 9'b011011001;
      9'b110011010: out = 9'b011011001; // overlap
      9'b110011011: out = 9'b011011010;
      9'b110011100: out = 9'b011011010; // overlap
      9'b110011101: out = 9'b011011010; // overlap
      9'b110011110: out = 9'b011011011;
      9'b110011111: out = 9'b011011011; // overlap
      9'b110100000: out = 9'b011011100;
      9'b110100001: out = 9'b011011100; // overlap
      9'b110100010: out = 9'b011011100; // overlap
      9'b110100011: out = 9'b011011101;
      9'b110100100: out = 9'b011011101; // overlap
      9'b110100101: out = 9'b011011110;
      9'b110100110: out = 9'b011011110; // overlap
      9'b110100111: out = 9'b011011110; // overlap
      9'b110101000: out = 9'b011011111;
      9'b110101001: out = 9'b011011111; // overlap
      9'b110101010: out = 9'b011100000;
      9'b110101011: out = 9'b011100000; // overlap
      9'b110101100: out = 9'b011100000; // overlap
      9'b110101101: out = 9'b011100001;
      9'b110101110: out = 9'b011100001; // overlap
      9'b110101111: out = 9'b011100010;
      9'b110110000: out = 9'b011100010; // overlap
      9'b110110001: out = 9'b011100010; // overlap
      9'b110110010: out = 9'b011100011;
      9'b110110011: out = 9'b011100011; // overlap
      9'b110110100: out = 9'b011100100;
      9'b110110101: out = 9'b011100100; // overlap
      9'b110110110: out = 9'b011100100; // overlap
      9'b110110111: out = 9'b011100101;
      9'b110111000: out = 9'b011100101; // overlap
      9'b110111001: out = 9'b011100101; // overlap
      9'b110111010: out = 9'b011100110;
      9'b110111011: out = 9'b011100110; // overlap
      9'b110111100: out = 9'b011100111;
      9'b110111101: out = 9'b011100111; // overlap
      9'b110111110: out = 9'b011100111; // overlap
      9'b110111111: out = 9'b011101000;
      9'b111000000: out = 9'b011101000; // overlap
      9'b111000001: out = 9'b011101001;
      9'b111000010: out = 9'b011101001; // overlap
      9'b111000011: out = 9'b011101001; // overlap
      9'b111000100: out = 9'b011101010;
      9'b111000101: out = 9'b011101010; // overlap
      9'b111000110: out = 9'b011101010; // overlap
      9'b111000111: out = 9'b011101011;
      9'b111001000: out = 9'b011101011; // overlap
      9'b111001001: out = 9'b011101100;
      9'b111001010: out = 9'b011101100; // overlap
      9'b111001011: out = 9'b011101100; // overlap
      9'b111001100: out = 9'b011101101;
      9'b111001101: out = 9'b011101101; // overlap
      9'b111001110: out = 9'b011101110;
      9'b111001111: out = 9'b011101110; // overlap
      9'b111010000: out = 9'b011101110; // overlap
      9'b111010001: out = 9'b011101111;
      9'b111010010: out = 9'b011101111; // overlap
      9'b111010011: out = 9'b011101111; // overlap
      9'b111010100: out = 9'b011110000;
      9'b111010101: out = 9'b011110000; // overlap
      9'b111010110: out = 9'b011110001;
      9'b111010111: out = 9'b011110001; // overlap
      9'b111011000: out = 9'b011110001; // overlap
      9'b111011001: out = 9'b011110010;
      9'b111011010: out = 9'b011110010; // overlap
      9'b111011011: out = 9'b011110010; // overlap
      9'b111011100: out = 9'b011110011;
      9'b111011101: out = 9'b011110011; // overlap
      9'b111011110: out = 9'b011110100;
      9'b111011111: out = 9'b011110100; // overlap
      9'b111100000: out = 9'b011110100; // overlap
      9'b111100001: out = 9'b011110101;
      9'b111100010: out = 9'b011110101; // overlap
      9'b111100011: out = 9'b011110101; // overlap
      9'b111100100: out = 9'b011110110;
      9'b111100101: out = 9'b011110110; // overlap
      9'b111100110: out = 9'b011110111;
      9'b111100111: out = 9'b011110111; // overlap
      9'b111101000: out = 9'b011110111; // overlap
      9'b111101001: out = 9'b011111000;
      9'b111101010: out = 9'b011111000; // overlap
      9'b111101011: out = 9'b011111000; // overlap
      9'b111101100: out = 9'b011111001;
      9'b111101101: out = 9'b011111001; // overlap
      9'b111101110: out = 9'b011111001; // overlap
      9'b111101111: out = 9'b011111010;
      9'b111110000: out = 9'b011111010; // overlap
      9'b111110001: out = 9'b011111011;
      9'b111110010: out = 9'b011111011; // overlap
      9'b111110011: out = 9'b011111011; // overlap
      9'b111110100: out = 9'b011111100;
      9'b111110101: out = 9'b011111100; // overlap
      9'b111110110: out = 9'b011111100; // overlap
      9'b111110111: out = 9'b011111101;
      9'b111111000: out = 9'b011111101; // overlap
      9'b111111001: out = 9'b011111101; // overlap
      9'b111111010: out = 9'b011111110;
      9'b111111011: out = 9'b011111110; // overlap
      9'b111111100: out = 9'b011111111;
      9'b111111101: out = 9'b011111111; // overlap
      9'b111111110: out = 9'b011111111; // overlap
      9'b111111111: out = 9'b100000000; // overlap + round
      default: out = 9'bxxxxxxxxx;
    endcase
  end
endmodule
