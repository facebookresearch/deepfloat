// Copyright (c) Facebook, Inc. and its affiliates. All Rights Reserved.
// All rights reserved.
//
// This source code is licensed under the license found in the
// LICENSE file in the root directory of this source tree.


module Pow2LUT_10x11
  (input [9:0] in,
   output logic [10:0] out);

  always_comb begin
    case (in)
      10'b0000000000: out = 11'b00000000000;
      10'b0000000001: out = 11'b00000000001;
      10'b0000000010: out = 11'b00000000011; // round
      10'b0000000011: out = 11'b00000000100;
      10'b0000000100: out = 11'b00000000110; // round
      10'b0000000101: out = 11'b00000000111; // round
      10'b0000000110: out = 11'b00000001000;
      10'b0000000111: out = 11'b00000001010; // round
      10'b0000001000: out = 11'b00000001011;
      10'b0000001001: out = 11'b00000001101; // round
      10'b0000001010: out = 11'b00000001110; // round
      10'b0000001011: out = 11'b00000001111;
      10'b0000001100: out = 11'b00000010001; // round
      10'b0000001101: out = 11'b00000010010;
      10'b0000001110: out = 11'b00000010100; // round
      10'b0000001111: out = 11'b00000010101; // round
      10'b0000010000: out = 11'b00000010110;
      10'b0000010001: out = 11'b00000011000; // round
      10'b0000010010: out = 11'b00000011001;
      10'b0000010011: out = 11'b00000011011; // round
      10'b0000010100: out = 11'b00000011100; // round
      10'b0000010101: out = 11'b00000011101;
      10'b0000010110: out = 11'b00000011111; // round
      10'b0000010111: out = 11'b00000100000;
      10'b0000011000: out = 11'b00000100010; // round
      10'b0000011001: out = 11'b00000100011; // round
      10'b0000011010: out = 11'b00000100100;
      10'b0000011011: out = 11'b00000100110; // round
      10'b0000011100: out = 11'b00000100111;
      10'b0000011101: out = 11'b00000101001; // round
      10'b0000011110: out = 11'b00000101010;
      10'b0000011111: out = 11'b00000101011;
      10'b0000100000: out = 11'b00000101101; // round
      10'b0000100001: out = 11'b00000101110;
      10'b0000100010: out = 11'b00000110000; // round
      10'b0000100011: out = 11'b00000110001;
      10'b0000100100: out = 11'b00000110011; // round
      10'b0000100101: out = 11'b00000110100; // round
      10'b0000100110: out = 11'b00000110101;
      10'b0000100111: out = 11'b00000110111; // round
      10'b0000101000: out = 11'b00000111000;
      10'b0000101001: out = 11'b00000111010; // round
      10'b0000101010: out = 11'b00000111011;
      10'b0000101011: out = 11'b00000111100;
      10'b0000101100: out = 11'b00000111110; // round
      10'b0000101101: out = 11'b00000111111;
      10'b0000101110: out = 11'b00001000001; // round
      10'b0000101111: out = 11'b00001000010;
      10'b0000110000: out = 11'b00001000100; // round
      10'b0000110001: out = 11'b00001000101;
      10'b0000110010: out = 11'b00001000111; // round
      10'b0000110011: out = 11'b00001001000; // round
      10'b0000110100: out = 11'b00001001001;
      10'b0000110101: out = 11'b00001001011; // round
      10'b0000110110: out = 11'b00001001100;
      10'b0000110111: out = 11'b00001001110; // round
      10'b0000111000: out = 11'b00001001111;
      10'b0000111001: out = 11'b00001010001; // round
      10'b0000111010: out = 11'b00001010010;
      10'b0000111011: out = 11'b00001010011;
      10'b0000111100: out = 11'b00001010101; // round
      10'b0000111101: out = 11'b00001010110;
      10'b0000111110: out = 11'b00001011000; // round
      10'b0000111111: out = 11'b00001011001;
      10'b0001000000: out = 11'b00001011011; // round
      10'b0001000001: out = 11'b00001011100;
      10'b0001000010: out = 11'b00001011110; // round
      10'b0001000011: out = 11'b00001011111;
      10'b0001000100: out = 11'b00001100000;
      10'b0001000101: out = 11'b00001100010; // round
      10'b0001000110: out = 11'b00001100011;
      10'b0001000111: out = 11'b00001100101; // round
      10'b0001001000: out = 11'b00001100110;
      10'b0001001001: out = 11'b00001101000; // round
      10'b0001001010: out = 11'b00001101001;
      10'b0001001011: out = 11'b00001101011; // round
      10'b0001001100: out = 11'b00001101100;
      10'b0001001101: out = 11'b00001101110; // round
      10'b0001001110: out = 11'b00001101111;
      10'b0001001111: out = 11'b00001110000;
      10'b0001010000: out = 11'b00001110010; // round
      10'b0001010001: out = 11'b00001110011;
      10'b0001010010: out = 11'b00001110101; // round
      10'b0001010011: out = 11'b00001110110;
      10'b0001010100: out = 11'b00001111000; // round
      10'b0001010101: out = 11'b00001111001;
      10'b0001010110: out = 11'b00001111011; // round
      10'b0001010111: out = 11'b00001111100;
      10'b0001011000: out = 11'b00001111110; // round
      10'b0001011001: out = 11'b00001111111;
      10'b0001011010: out = 11'b00010000001; // round
      10'b0001011011: out = 11'b00010000010;
      10'b0001011100: out = 11'b00010000100; // round
      10'b0001011101: out = 11'b00010000101;
      10'b0001011110: out = 11'b00010000111; // round
      10'b0001011111: out = 11'b00010001000;
      10'b0001100000: out = 11'b00010001010; // round
      10'b0001100001: out = 11'b00010001011; // round
      10'b0001100010: out = 11'b00010001100;
      10'b0001100011: out = 11'b00010001110; // round
      10'b0001100100: out = 11'b00010001111;
      10'b0001100101: out = 11'b00010010001; // round
      10'b0001100110: out = 11'b00010010010;
      10'b0001100111: out = 11'b00010010100; // round
      10'b0001101000: out = 11'b00010010101;
      10'b0001101001: out = 11'b00010010111; // round
      10'b0001101010: out = 11'b00010011000;
      10'b0001101011: out = 11'b00010011010; // round
      10'b0001101100: out = 11'b00010011011;
      10'b0001101101: out = 11'b00010011101; // round
      10'b0001101110: out = 11'b00010011110;
      10'b0001101111: out = 11'b00010100000; // round
      10'b0001110000: out = 11'b00010100001;
      10'b0001110001: out = 11'b00010100011; // round
      10'b0001110010: out = 11'b00010100100;
      10'b0001110011: out = 11'b00010100110; // round
      10'b0001110100: out = 11'b00010100111;
      10'b0001110101: out = 11'b00010101001; // round
      10'b0001110110: out = 11'b00010101010;
      10'b0001110111: out = 11'b00010101100; // round
      10'b0001111000: out = 11'b00010101101;
      10'b0001111001: out = 11'b00010101111; // round
      10'b0001111010: out = 11'b00010110000;
      10'b0001111011: out = 11'b00010110010; // round
      10'b0001111100: out = 11'b00010110011;
      10'b0001111101: out = 11'b00010110101; // round
      10'b0001111110: out = 11'b00010110110;
      10'b0001111111: out = 11'b00010111000; // round
      10'b0010000000: out = 11'b00010111001;
      10'b0010000001: out = 11'b00010111011; // round
      10'b0010000010: out = 11'b00010111100;
      10'b0010000011: out = 11'b00010111110; // round
      10'b0010000100: out = 11'b00010111111;
      10'b0010000101: out = 11'b00011000001; // round
      10'b0010000110: out = 11'b00011000010;
      10'b0010000111: out = 11'b00011000100; // round
      10'b0010001000: out = 11'b00011000101;
      10'b0010001001: out = 11'b00011000111;
      10'b0010001010: out = 11'b00011001001; // round
      10'b0010001011: out = 11'b00011001010;
      10'b0010001100: out = 11'b00011001100; // round
      10'b0010001101: out = 11'b00011001101;
      10'b0010001110: out = 11'b00011001111; // round
      10'b0010001111: out = 11'b00011010000;
      10'b0010010000: out = 11'b00011010010; // round
      10'b0010010001: out = 11'b00011010011;
      10'b0010010010: out = 11'b00011010101; // round
      10'b0010010011: out = 11'b00011010110;
      10'b0010010100: out = 11'b00011011000; // round
      10'b0010010101: out = 11'b00011011001;
      10'b0010010110: out = 11'b00011011011; // round
      10'b0010010111: out = 11'b00011011100;
      10'b0010011000: out = 11'b00011011110; // round
      10'b0010011001: out = 11'b00011011111;
      10'b0010011010: out = 11'b00011100001;
      10'b0010011011: out = 11'b00011100011; // round
      10'b0010011100: out = 11'b00011100100;
      10'b0010011101: out = 11'b00011100110; // round
      10'b0010011110: out = 11'b00011100111;
      10'b0010011111: out = 11'b00011101001; // round
      10'b0010100000: out = 11'b00011101010;
      10'b0010100001: out = 11'b00011101100; // round
      10'b0010100010: out = 11'b00011101101;
      10'b0010100011: out = 11'b00011101111; // round
      10'b0010100100: out = 11'b00011110000;
      10'b0010100101: out = 11'b00011110010;
      10'b0010100110: out = 11'b00011110100; // round
      10'b0010100111: out = 11'b00011110101;
      10'b0010101000: out = 11'b00011110111; // round
      10'b0010101001: out = 11'b00011111000;
      10'b0010101010: out = 11'b00011111010; // round
      10'b0010101011: out = 11'b00011111011;
      10'b0010101100: out = 11'b00011111101; // round
      10'b0010101101: out = 11'b00011111110;
      10'b0010101110: out = 11'b00100000000; // round
      10'b0010101111: out = 11'b00100000010; // round
      10'b0010110000: out = 11'b00100000011;
      10'b0010110001: out = 11'b00100000101; // round
      10'b0010110010: out = 11'b00100000110;
      10'b0010110011: out = 11'b00100001000; // round
      10'b0010110100: out = 11'b00100001001;
      10'b0010110101: out = 11'b00100001011; // round
      10'b0010110110: out = 11'b00100001101; // round
      10'b0010110111: out = 11'b00100001110;
      10'b0010111000: out = 11'b00100010000; // round
      10'b0010111001: out = 11'b00100010001;
      10'b0010111010: out = 11'b00100010011; // round
      10'b0010111011: out = 11'b00100010100;
      10'b0010111100: out = 11'b00100010110; // round
      10'b0010111101: out = 11'b00100011000; // round
      10'b0010111110: out = 11'b00100011001;
      10'b0010111111: out = 11'b00100011011; // round
      10'b0011000000: out = 11'b00100011100;
      10'b0011000001: out = 11'b00100011110; // round
      10'b0011000010: out = 11'b00100011111;
      10'b0011000011: out = 11'b00100100001; // round
      10'b0011000100: out = 11'b00100100011; // round
      10'b0011000101: out = 11'b00100100100;
      10'b0011000110: out = 11'b00100100110; // round
      10'b0011000111: out = 11'b00100100111;
      10'b0011001000: out = 11'b00100101001; // round
      10'b0011001001: out = 11'b00100101010;
      10'b0011001010: out = 11'b00100101100;
      10'b0011001011: out = 11'b00100101110; // round
      10'b0011001100: out = 11'b00100101111;
      10'b0011001101: out = 11'b00100110001; // round
      10'b0011001110: out = 11'b00100110010;
      10'b0011001111: out = 11'b00100110100;
      10'b0011010000: out = 11'b00100110110; // round
      10'b0011010001: out = 11'b00100110111;
      10'b0011010010: out = 11'b00100111001; // round
      10'b0011010011: out = 11'b00100111010;
      10'b0011010100: out = 11'b00100111100;
      10'b0011010101: out = 11'b00100111110; // round
      10'b0011010110: out = 11'b00100111111;
      10'b0011010111: out = 11'b00101000001; // round
      10'b0011011000: out = 11'b00101000010;
      10'b0011011001: out = 11'b00101000100;
      10'b0011011010: out = 11'b00101000110; // round
      10'b0011011011: out = 11'b00101000111;
      10'b0011011100: out = 11'b00101001001; // round
      10'b0011011101: out = 11'b00101001010;
      10'b0011011110: out = 11'b00101001100;
      10'b0011011111: out = 11'b00101001110; // round
      10'b0011100000: out = 11'b00101001111;
      10'b0011100001: out = 11'b00101010001; // round
      10'b0011100010: out = 11'b00101010011; // round
      10'b0011100011: out = 11'b00101010100;
      10'b0011100100: out = 11'b00101010110; // round
      10'b0011100101: out = 11'b00101010111;
      10'b0011100110: out = 11'b00101011001;
      10'b0011100111: out = 11'b00101011011; // round
      10'b0011101000: out = 11'b00101011100;
      10'b0011101001: out = 11'b00101011110; // round
      10'b0011101010: out = 11'b00101011111;
      10'b0011101011: out = 11'b00101100001;
      10'b0011101100: out = 11'b00101100011; // round
      10'b0011101101: out = 11'b00101100100;
      10'b0011101110: out = 11'b00101100110;
      10'b0011101111: out = 11'b00101101000; // round
      10'b0011110000: out = 11'b00101101001;
      10'b0011110001: out = 11'b00101101011; // round
      10'b0011110010: out = 11'b00101101101; // round
      10'b0011110011: out = 11'b00101101110;
      10'b0011110100: out = 11'b00101110000; // round
      10'b0011110101: out = 11'b00101110001;
      10'b0011110110: out = 11'b00101110011;
      10'b0011110111: out = 11'b00101110101; // round
      10'b0011111000: out = 11'b00101110110;
      10'b0011111001: out = 11'b00101111000; // round
      10'b0011111010: out = 11'b00101111010; // round
      10'b0011111011: out = 11'b00101111011;
      10'b0011111100: out = 11'b00101111101; // round
      10'b0011111101: out = 11'b00101111111; // round
      10'b0011111110: out = 11'b00110000000;
      10'b0011111111: out = 11'b00110000010; // round
      10'b0100000000: out = 11'b00110000011;
      10'b0100000001: out = 11'b00110000101;
      10'b0100000010: out = 11'b00110000111; // round
      10'b0100000011: out = 11'b00110001000;
      10'b0100000100: out = 11'b00110001010;
      10'b0100000101: out = 11'b00110001100; // round
      10'b0100000110: out = 11'b00110001101;
      10'b0100000111: out = 11'b00110001111;
      10'b0100001000: out = 11'b00110010001; // round
      10'b0100001001: out = 11'b00110010010;
      10'b0100001010: out = 11'b00110010100;
      10'b0100001011: out = 11'b00110010110; // round
      10'b0100001100: out = 11'b00110010111;
      10'b0100001101: out = 11'b00110011001;
      10'b0100001110: out = 11'b00110011011; // round
      10'b0100001111: out = 11'b00110011100;
      10'b0100010000: out = 11'b00110011110;
      10'b0100010001: out = 11'b00110100000; // round
      10'b0100010010: out = 11'b00110100001;
      10'b0100010011: out = 11'b00110100011;
      10'b0100010100: out = 11'b00110100101; // round
      10'b0100010101: out = 11'b00110100110;
      10'b0100010110: out = 11'b00110101000;
      10'b0100010111: out = 11'b00110101010; // round
      10'b0100011000: out = 11'b00110101011;
      10'b0100011001: out = 11'b00110101101;
      10'b0100011010: out = 11'b00110101111; // round
      10'b0100011011: out = 11'b00110110000;
      10'b0100011100: out = 11'b00110110010;
      10'b0100011101: out = 11'b00110110100; // round
      10'b0100011110: out = 11'b00110110101;
      10'b0100011111: out = 11'b00110110111;
      10'b0100100000: out = 11'b00110111001; // round
      10'b0100100001: out = 11'b00110111011; // round
      10'b0100100010: out = 11'b00110111100;
      10'b0100100011: out = 11'b00110111110; // round
      10'b0100100100: out = 11'b00111000000; // round
      10'b0100100101: out = 11'b00111000001;
      10'b0100100110: out = 11'b00111000011; // round
      10'b0100100111: out = 11'b00111000101; // round
      10'b0100101000: out = 11'b00111000110;
      10'b0100101001: out = 11'b00111001000;
      10'b0100101010: out = 11'b00111001010; // round
      10'b0100101011: out = 11'b00111001011;
      10'b0100101100: out = 11'b00111001101;
      10'b0100101101: out = 11'b00111001111; // round
      10'b0100101110: out = 11'b00111010001; // round
      10'b0100101111: out = 11'b00111010010;
      10'b0100110000: out = 11'b00111010100; // round
      10'b0100110001: out = 11'b00111010110; // round
      10'b0100110010: out = 11'b00111010111;
      10'b0100110011: out = 11'b00111011001;
      10'b0100110100: out = 11'b00111011011; // round
      10'b0100110101: out = 11'b00111011100;
      10'b0100110110: out = 11'b00111011110;
      10'b0100110111: out = 11'b00111100000; // round
      10'b0100111000: out = 11'b00111100010; // round
      10'b0100111001: out = 11'b00111100011;
      10'b0100111010: out = 11'b00111100101;
      10'b0100111011: out = 11'b00111100111; // round
      10'b0100111100: out = 11'b00111101000;
      10'b0100111101: out = 11'b00111101010;
      10'b0100111110: out = 11'b00111101100; // round
      10'b0100111111: out = 11'b00111101110; // round
      10'b0101000000: out = 11'b00111101111;
      10'b0101000001: out = 11'b00111110001;
      10'b0101000010: out = 11'b00111110011; // round
      10'b0101000011: out = 11'b00111110100;
      10'b0101000100: out = 11'b00111110110;
      10'b0101000101: out = 11'b00111111000; // round
      10'b0101000110: out = 11'b00111111010; // round
      10'b0101000111: out = 11'b00111111011;
      10'b0101001000: out = 11'b00111111101;
      10'b0101001001: out = 11'b00111111111; // round
      10'b0101001010: out = 11'b01000000001; // round
      10'b0101001011: out = 11'b01000000010;
      10'b0101001100: out = 11'b01000000100;
      10'b0101001101: out = 11'b01000000110; // round
      10'b0101001110: out = 11'b01000001000; // round
      10'b0101001111: out = 11'b01000001001;
      10'b0101010000: out = 11'b01000001011;
      10'b0101010001: out = 11'b01000001101; // round
      10'b0101010010: out = 11'b01000001111; // round
      10'b0101010011: out = 11'b01000010000;
      10'b0101010100: out = 11'b01000010010; // round
      10'b0101010101: out = 11'b01000010100; // round
      10'b0101010110: out = 11'b01000010101;
      10'b0101010111: out = 11'b01000010111;
      10'b0101011000: out = 11'b01000011001; // round
      10'b0101011001: out = 11'b01000011011; // round
      10'b0101011010: out = 11'b01000011100;
      10'b0101011011: out = 11'b01000011110;
      10'b0101011100: out = 11'b01000100000; // round
      10'b0101011101: out = 11'b01000100010; // round
      10'b0101011110: out = 11'b01000100100; // round
      10'b0101011111: out = 11'b01000100101;
      10'b0101100000: out = 11'b01000100111;
      10'b0101100001: out = 11'b01000101001; // round
      10'b0101100010: out = 11'b01000101011; // round
      10'b0101100011: out = 11'b01000101100;
      10'b0101100100: out = 11'b01000101110;
      10'b0101100101: out = 11'b01000110000; // round
      10'b0101100110: out = 11'b01000110010; // round
      10'b0101100111: out = 11'b01000110011;
      10'b0101101000: out = 11'b01000110101;
      10'b0101101001: out = 11'b01000110111; // round
      10'b0101101010: out = 11'b01000111001; // round
      10'b0101101011: out = 11'b01000111010;
      10'b0101101100: out = 11'b01000111100;
      10'b0101101101: out = 11'b01000111110; // round
      10'b0101101110: out = 11'b01001000000; // round
      10'b0101101111: out = 11'b01001000010; // round
      10'b0101110000: out = 11'b01001000011;
      10'b0101110001: out = 11'b01001000101;
      10'b0101110010: out = 11'b01001000111; // round
      10'b0101110011: out = 11'b01001001001; // round
      10'b0101110100: out = 11'b01001001010;
      10'b0101110101: out = 11'b01001001100;
      10'b0101110110: out = 11'b01001001110;
      10'b0101110111: out = 11'b01001010000; // round
      10'b0101111000: out = 11'b01001010010; // round
      10'b0101111001: out = 11'b01001010011;
      10'b0101111010: out = 11'b01001010101;
      10'b0101111011: out = 11'b01001010111; // round
      10'b0101111100: out = 11'b01001011001; // round
      10'b0101111101: out = 11'b01001011011; // round
      10'b0101111110: out = 11'b01001011100;
      10'b0101111111: out = 11'b01001011110;
      10'b0110000000: out = 11'b01001100000; // round
      10'b0110000001: out = 11'b01001100010; // round
      10'b0110000010: out = 11'b01001100100; // round
      10'b0110000011: out = 11'b01001100101;
      10'b0110000100: out = 11'b01001100111;
      10'b0110000101: out = 11'b01001101001; // round
      10'b0110000110: out = 11'b01001101011; // round
      10'b0110000111: out = 11'b01001101101; // round
      10'b0110001000: out = 11'b01001101110;
      10'b0110001001: out = 11'b01001110000;
      10'b0110001010: out = 11'b01001110010; // round
      10'b0110001011: out = 11'b01001110100; // round
      10'b0110001100: out = 11'b01001110110; // round
      10'b0110001101: out = 11'b01001110111;
      10'b0110001110: out = 11'b01001111001;
      10'b0110001111: out = 11'b01001111011;
      10'b0110010000: out = 11'b01001111101; // round
      10'b0110010001: out = 11'b01001111111; // round
      10'b0110010010: out = 11'b01010000000;
      10'b0110010011: out = 11'b01010000010;
      10'b0110010100: out = 11'b01010000100;
      10'b0110010101: out = 11'b01010000110; // round
      10'b0110010110: out = 11'b01010001000; // round
      10'b0110010111: out = 11'b01010001010; // round
      10'b0110011000: out = 11'b01010001011;
      10'b0110011001: out = 11'b01010001101;
      10'b0110011010: out = 11'b01010001111;
      10'b0110011011: out = 11'b01010010001; // round
      10'b0110011100: out = 11'b01010010011; // round
      10'b0110011101: out = 11'b01010010101; // round
      10'b0110011110: out = 11'b01010010110;
      10'b0110011111: out = 11'b01010011000;
      10'b0110100000: out = 11'b01010011010;
      10'b0110100001: out = 11'b01010011100; // round
      10'b0110100010: out = 11'b01010011110; // round
      10'b0110100011: out = 11'b01010100000; // round
      10'b0110100100: out = 11'b01010100001;
      10'b0110100101: out = 11'b01010100011;
      10'b0110100110: out = 11'b01010100101;
      10'b0110100111: out = 11'b01010100111; // round
      10'b0110101000: out = 11'b01010101001; // round
      10'b0110101001: out = 11'b01010101011; // round
      10'b0110101010: out = 11'b01010101101; // round
      10'b0110101011: out = 11'b01010101110;
      10'b0110101100: out = 11'b01010110000;
      10'b0110101101: out = 11'b01010110010;
      10'b0110101110: out = 11'b01010110100; // round
      10'b0110101111: out = 11'b01010110110; // round
      10'b0110110000: out = 11'b01010111000; // round
      10'b0110110001: out = 11'b01010111001;
      10'b0110110010: out = 11'b01010111011;
      10'b0110110011: out = 11'b01010111101;
      10'b0110110100: out = 11'b01010111111;
      10'b0110110101: out = 11'b01011000001; // round
      10'b0110110110: out = 11'b01011000011; // round
      10'b0110110111: out = 11'b01011000101; // round
      10'b0110111000: out = 11'b01011000111; // round
      10'b0110111001: out = 11'b01011001000;
      10'b0110111010: out = 11'b01011001010;
      10'b0110111011: out = 11'b01011001100;
      10'b0110111100: out = 11'b01011001110;
      10'b0110111101: out = 11'b01011010000; // round
      10'b0110111110: out = 11'b01011010010; // round
      10'b0110111111: out = 11'b01011010100; // round
      10'b0111000000: out = 11'b01011010110; // round
      10'b0111000001: out = 11'b01011010111;
      10'b0111000010: out = 11'b01011011001;
      10'b0111000011: out = 11'b01011011011;
      10'b0111000100: out = 11'b01011011101;
      10'b0111000101: out = 11'b01011011111; // round
      10'b0111000110: out = 11'b01011100001; // round
      10'b0111000111: out = 11'b01011100011; // round
      10'b0111001000: out = 11'b01011100101; // round
      10'b0111001001: out = 11'b01011100110;
      10'b0111001010: out = 11'b01011101000;
      10'b0111001011: out = 11'b01011101010;
      10'b0111001100: out = 11'b01011101100;
      10'b0111001101: out = 11'b01011101110;
      10'b0111001110: out = 11'b01011110000; // round
      10'b0111001111: out = 11'b01011110010; // round
      10'b0111010000: out = 11'b01011110100; // round
      10'b0111010001: out = 11'b01011110110; // round
      10'b0111010010: out = 11'b01011111000; // round
      10'b0111010011: out = 11'b01011111001;
      10'b0111010100: out = 11'b01011111011;
      10'b0111010101: out = 11'b01011111101;
      10'b0111010110: out = 11'b01011111111;
      10'b0111010111: out = 11'b01100000001;
      10'b0111011000: out = 11'b01100000011; // round
      10'b0111011001: out = 11'b01100000101; // round
      10'b0111011010: out = 11'b01100000111; // round
      10'b0111011011: out = 11'b01100001001; // round
      10'b0111011100: out = 11'b01100001011; // round
      10'b0111011101: out = 11'b01100001100;
      10'b0111011110: out = 11'b01100001110;
      10'b0111011111: out = 11'b01100010000;
      10'b0111100000: out = 11'b01100010010;
      10'b0111100001: out = 11'b01100010100;
      10'b0111100010: out = 11'b01100010110;
      10'b0111100011: out = 11'b01100011000;
      10'b0111100100: out = 11'b01100011010; // round
      10'b0111100101: out = 11'b01100011100; // round
      10'b0111100110: out = 11'b01100011110; // round
      10'b0111100111: out = 11'b01100100000; // round
      10'b0111101000: out = 11'b01100100010; // round
      10'b0111101001: out = 11'b01100100100; // round
      10'b0111101010: out = 11'b01100100101;
      10'b0111101011: out = 11'b01100100111;
      10'b0111101100: out = 11'b01100101001;
      10'b0111101101: out = 11'b01100101011;
      10'b0111101110: out = 11'b01100101101;
      10'b0111101111: out = 11'b01100101111;
      10'b0111110000: out = 11'b01100110001;
      10'b0111110001: out = 11'b01100110011;
      10'b0111110010: out = 11'b01100110101; // round
      10'b0111110011: out = 11'b01100110111; // round
      10'b0111110100: out = 11'b01100111001; // round
      10'b0111110101: out = 11'b01100111011; // round
      10'b0111110110: out = 11'b01100111101; // round
      10'b0111110111: out = 11'b01100111111; // round
      10'b0111111000: out = 11'b01101000001; // round
      10'b0111111001: out = 11'b01101000011; // round
      10'b0111111010: out = 11'b01101000101; // round
      10'b0111111011: out = 11'b01101000111; // round
      10'b0111111100: out = 11'b01101001000;
      10'b0111111101: out = 11'b01101001010;
      10'b0111111110: out = 11'b01101001100;
      10'b0111111111: out = 11'b01101001110;
      10'b1000000000: out = 11'b01101010000;
      10'b1000000001: out = 11'b01101010010;
      10'b1000000010: out = 11'b01101010100;
      10'b1000000011: out = 11'b01101010110;
      10'b1000000100: out = 11'b01101011000;
      10'b1000000101: out = 11'b01101011010;
      10'b1000000110: out = 11'b01101011100;
      10'b1000000111: out = 11'b01101011110;
      10'b1000001000: out = 11'b01101100000;
      10'b1000001001: out = 11'b01101100010;
      10'b1000001010: out = 11'b01101100100; // round
      10'b1000001011: out = 11'b01101100110; // round
      10'b1000001100: out = 11'b01101101000; // round
      10'b1000001101: out = 11'b01101101010; // round
      10'b1000001110: out = 11'b01101101100; // round
      10'b1000001111: out = 11'b01101101110; // round
      10'b1000010000: out = 11'b01101110000; // round
      10'b1000010001: out = 11'b01101110010; // round
      10'b1000010010: out = 11'b01101110100; // round
      10'b1000010011: out = 11'b01101110110; // round
      10'b1000010100: out = 11'b01101111000; // round
      10'b1000010101: out = 11'b01101111010; // round
      10'b1000010110: out = 11'b01101111100; // round
      10'b1000010111: out = 11'b01101111110; // round
      10'b1000011000: out = 11'b01110000000; // round
      10'b1000011001: out = 11'b01110000010; // round
      10'b1000011010: out = 11'b01110000100; // round
      10'b1000011011: out = 11'b01110000110; // round
      10'b1000011100: out = 11'b01110001000; // round
      10'b1000011101: out = 11'b01110001010; // round
      10'b1000011110: out = 11'b01110001100; // round
      10'b1000011111: out = 11'b01110001110; // round
      10'b1000100000: out = 11'b01110010000; // round
      10'b1000100001: out = 11'b01110010010; // round
      10'b1000100010: out = 11'b01110010100; // round
      10'b1000100011: out = 11'b01110010110; // round
      10'b1000100100: out = 11'b01110011000; // round
      10'b1000100101: out = 11'b01110011010; // round
      10'b1000100110: out = 11'b01110011100; // round
      10'b1000100111: out = 11'b01110011110; // round
      10'b1000101000: out = 11'b01110100000; // round
      10'b1000101001: out = 11'b01110100010; // round
      10'b1000101010: out = 11'b01110100100; // round
      10'b1000101011: out = 11'b01110100110; // round
      10'b1000101100: out = 11'b01110101000; // round
      10'b1000101101: out = 11'b01110101010; // round
      10'b1000101110: out = 11'b01110101100; // round
      10'b1000101111: out = 11'b01110101110; // round
      10'b1000110000: out = 11'b01110110000; // round
      10'b1000110001: out = 11'b01110110010; // round
      10'b1000110010: out = 11'b01110110100;
      10'b1000110011: out = 11'b01110110110;
      10'b1000110100: out = 11'b01110111000;
      10'b1000110101: out = 11'b01110111010;
      10'b1000110110: out = 11'b01110111100;
      10'b1000110111: out = 11'b01110111110;
      10'b1000111000: out = 11'b01111000000;
      10'b1000111001: out = 11'b01111000010;
      10'b1000111010: out = 11'b01111000100;
      10'b1000111011: out = 11'b01111000110;
      10'b1000111100: out = 11'b01111001000;
      10'b1000111101: out = 11'b01111001010;
      10'b1000111110: out = 11'b01111001100;
      10'b1000111111: out = 11'b01111001110;
      10'b1001000000: out = 11'b01111010001; // round
      10'b1001000001: out = 11'b01111010011; // round
      10'b1001000010: out = 11'b01111010101; // round
      10'b1001000011: out = 11'b01111010111; // round
      10'b1001000100: out = 11'b01111011001; // round
      10'b1001000101: out = 11'b01111011011; // round
      10'b1001000110: out = 11'b01111011101; // round
      10'b1001000111: out = 11'b01111011111; // round
      10'b1001001000: out = 11'b01111100001; // round
      10'b1001001001: out = 11'b01111100011;
      10'b1001001010: out = 11'b01111100101;
      10'b1001001011: out = 11'b01111100111;
      10'b1001001100: out = 11'b01111101001;
      10'b1001001101: out = 11'b01111101011;
      10'b1001001110: out = 11'b01111101101;
      10'b1001001111: out = 11'b01111101111;
      10'b1001010000: out = 11'b01111110001;
      10'b1001010001: out = 11'b01111110100; // round
      10'b1001010010: out = 11'b01111110110; // round
      10'b1001010011: out = 11'b01111111000; // round
      10'b1001010100: out = 11'b01111111010; // round
      10'b1001010101: out = 11'b01111111100; // round
      10'b1001010110: out = 11'b01111111110; // round
      10'b1001010111: out = 11'b10000000000; // round
      10'b1001011000: out = 11'b10000000010;
      10'b1001011001: out = 11'b10000000100;
      10'b1001011010: out = 11'b10000000110;
      10'b1001011011: out = 11'b10000001000;
      10'b1001011100: out = 11'b10000001010;
      10'b1001011101: out = 11'b10000001100;
      10'b1001011110: out = 11'b10000001111; // round
      10'b1001011111: out = 11'b10000010001; // round
      10'b1001100000: out = 11'b10000010011; // round
      10'b1001100001: out = 11'b10000010101; // round
      10'b1001100010: out = 11'b10000010111; // round
      10'b1001100011: out = 11'b10000011001;
      10'b1001100100: out = 11'b10000011011;
      10'b1001100101: out = 11'b10000011101;
      10'b1001100110: out = 11'b10000011111;
      10'b1001100111: out = 11'b10000100001;
      10'b1001101000: out = 11'b10000100100; // round
      10'b1001101001: out = 11'b10000100110; // round
      10'b1001101010: out = 11'b10000101000; // round
      10'b1001101011: out = 11'b10000101010; // round
      10'b1001101100: out = 11'b10000101100; // round
      10'b1001101101: out = 11'b10000101110;
      10'b1001101110: out = 11'b10000110000;
      10'b1001101111: out = 11'b10000110010;
      10'b1001110000: out = 11'b10000110100;
      10'b1001110001: out = 11'b10000110111; // round
      10'b1001110010: out = 11'b10000111001; // round
      10'b1001110011: out = 11'b10000111011; // round
      10'b1001110100: out = 11'b10000111101; // round
      10'b1001110101: out = 11'b10000111111;
      10'b1001110110: out = 11'b10001000001;
      10'b1001110111: out = 11'b10001000011;
      10'b1001111000: out = 11'b10001000101;
      10'b1001111001: out = 11'b10001001000; // round
      10'b1001111010: out = 11'b10001001010; // round
      10'b1001111011: out = 11'b10001001100; // round
      10'b1001111100: out = 11'b10001001110; // round
      10'b1001111101: out = 11'b10001010000;
      10'b1001111110: out = 11'b10001010010;
      10'b1001111111: out = 11'b10001010100;
      10'b1010000000: out = 11'b10001010110;
      10'b1010000001: out = 11'b10001011001; // round
      10'b1010000010: out = 11'b10001011011; // round
      10'b1010000011: out = 11'b10001011101; // round
      10'b1010000100: out = 11'b10001011111;
      10'b1010000101: out = 11'b10001100001;
      10'b1010000110: out = 11'b10001100011;
      10'b1010000111: out = 11'b10001100101;
      10'b1010001000: out = 11'b10001101000; // round
      10'b1010001001: out = 11'b10001101010; // round
      10'b1010001010: out = 11'b10001101100; // round
      10'b1010001011: out = 11'b10001101110;
      10'b1010001100: out = 11'b10001110000;
      10'b1010001101: out = 11'b10001110010;
      10'b1010001110: out = 11'b10001110101; // round
      10'b1010001111: out = 11'b10001110111; // round
      10'b1010010000: out = 11'b10001111001; // round
      10'b1010010001: out = 11'b10001111011;
      10'b1010010010: out = 11'b10001111101;
      10'b1010010011: out = 11'b10001111111;
      10'b1010010100: out = 11'b10010000001;
      10'b1010010101: out = 11'b10010000100; // round
      10'b1010010110: out = 11'b10010000110; // round
      10'b1010010111: out = 11'b10010001000;
      10'b1010011000: out = 11'b10010001010;
      10'b1010011001: out = 11'b10010001100;
      10'b1010011010: out = 11'b10010001111; // round
      10'b1010011011: out = 11'b10010010001; // round
      10'b1010011100: out = 11'b10010010011; // round
      10'b1010011101: out = 11'b10010010101;
      10'b1010011110: out = 11'b10010010111;
      10'b1010011111: out = 11'b10010011001;
      10'b1010100000: out = 11'b10010011100; // round
      10'b1010100001: out = 11'b10010011110; // round
      10'b1010100010: out = 11'b10010100000; // round
      10'b1010100011: out = 11'b10010100010;
      10'b1010100100: out = 11'b10010100100;
      10'b1010100101: out = 11'b10010100111; // round
      10'b1010100110: out = 11'b10010101001; // round
      10'b1010100111: out = 11'b10010101011; // round
      10'b1010101000: out = 11'b10010101101;
      10'b1010101001: out = 11'b10010101111;
      10'b1010101010: out = 11'b10010110010; // round
      10'b1010101011: out = 11'b10010110100; // round
      10'b1010101100: out = 11'b10010110110; // round
      10'b1010101101: out = 11'b10010111000;
      10'b1010101110: out = 11'b10010111010;
      10'b1010101111: out = 11'b10010111101; // round
      10'b1010110000: out = 11'b10010111111; // round
      10'b1010110001: out = 11'b10011000001; // round
      10'b1010110010: out = 11'b10011000011;
      10'b1010110011: out = 11'b10011000101;
      10'b1010110100: out = 11'b10011001000; // round
      10'b1010110101: out = 11'b10011001010; // round
      10'b1010110110: out = 11'b10011001100;
      10'b1010110111: out = 11'b10011001110;
      10'b1010111000: out = 11'b10011010000;
      10'b1010111001: out = 11'b10011010011; // round
      10'b1010111010: out = 11'b10011010101; // round
      10'b1010111011: out = 11'b10011010111;
      10'b1010111100: out = 11'b10011011001;
      10'b1010111101: out = 11'b10011011100; // round
      10'b1010111110: out = 11'b10011011110; // round
      10'b1010111111: out = 11'b10011100000;
      10'b1011000000: out = 11'b10011100010;
      10'b1011000001: out = 11'b10011100101; // round
      10'b1011000010: out = 11'b10011100111; // round
      10'b1011000011: out = 11'b10011101001; // round
      10'b1011000100: out = 11'b10011101011;
      10'b1011000101: out = 11'b10011101101;
      10'b1011000110: out = 11'b10011110000; // round
      10'b1011000111: out = 11'b10011110010; // round
      10'b1011001000: out = 11'b10011110100;
      10'b1011001001: out = 11'b10011110110;
      10'b1011001010: out = 11'b10011111001; // round
      10'b1011001011: out = 11'b10011111011; // round
      10'b1011001100: out = 11'b10011111101;
      10'b1011001101: out = 11'b10011111111;
      10'b1011001110: out = 11'b10100000010; // round
      10'b1011001111: out = 11'b10100000100; // round
      10'b1011010000: out = 11'b10100000110;
      10'b1011010001: out = 11'b10100001000;
      10'b1011010010: out = 11'b10100001011; // round
      10'b1011010011: out = 11'b10100001101; // round
      10'b1011010100: out = 11'b10100001111;
      10'b1011010101: out = 11'b10100010010; // round
      10'b1011010110: out = 11'b10100010100; // round
      10'b1011010111: out = 11'b10100010110;
      10'b1011011000: out = 11'b10100011000;
      10'b1011011001: out = 11'b10100011011; // round
      10'b1011011010: out = 11'b10100011101; // round
      10'b1011011011: out = 11'b10100011111;
      10'b1011011100: out = 11'b10100100001;
      10'b1011011101: out = 11'b10100100100; // round
      10'b1011011110: out = 11'b10100100110; // round
      10'b1011011111: out = 11'b10100101000;
      10'b1011100000: out = 11'b10100101011; // round
      10'b1011100001: out = 11'b10100101101; // round
      10'b1011100010: out = 11'b10100101111;
      10'b1011100011: out = 11'b10100110001;
      10'b1011100100: out = 11'b10100110100; // round
      10'b1011100101: out = 11'b10100110110; // round
      10'b1011100110: out = 11'b10100111000;
      10'b1011100111: out = 11'b10100111011; // round
      10'b1011101000: out = 11'b10100111101; // round
      10'b1011101001: out = 11'b10100111111;
      10'b1011101010: out = 11'b10101000001;
      10'b1011101011: out = 11'b10101000100; // round
      10'b1011101100: out = 11'b10101000110; // round
      10'b1011101101: out = 11'b10101001000;
      10'b1011101110: out = 11'b10101001011; // round
      10'b1011101111: out = 11'b10101001101; // round
      10'b1011110000: out = 11'b10101001111;
      10'b1011110001: out = 11'b10101010010; // round
      10'b1011110010: out = 11'b10101010100; // round
      10'b1011110011: out = 11'b10101010110;
      10'b1011110100: out = 11'b10101011000;
      10'b1011110101: out = 11'b10101011011; // round
      10'b1011110110: out = 11'b10101011101;
      10'b1011110111: out = 11'b10101011111;
      10'b1011111000: out = 11'b10101100010; // round
      10'b1011111001: out = 11'b10101100100;
      10'b1011111010: out = 11'b10101100110;
      10'b1011111011: out = 11'b10101101001; // round
      10'b1011111100: out = 11'b10101101011; // round
      10'b1011111101: out = 11'b10101101101;
      10'b1011111110: out = 11'b10101110000; // round
      10'b1011111111: out = 11'b10101110010; // round
      10'b1100000000: out = 11'b10101110100;
      10'b1100000001: out = 11'b10101110111; // round
      10'b1100000010: out = 11'b10101111001; // round
      10'b1100000011: out = 11'b10101111011;
      10'b1100000100: out = 11'b10101111110; // round
      10'b1100000101: out = 11'b10110000000; // round
      10'b1100000110: out = 11'b10110000010;
      10'b1100000111: out = 11'b10110000101; // round
      10'b1100001000: out = 11'b10110000111;
      10'b1100001001: out = 11'b10110001001;
      10'b1100001010: out = 11'b10110001100; // round
      10'b1100001011: out = 11'b10110001110;
      10'b1100001100: out = 11'b10110010000;
      10'b1100001101: out = 11'b10110010011; // round
      10'b1100001110: out = 11'b10110010101;
      10'b1100001111: out = 11'b10110010111;
      10'b1100010000: out = 11'b10110011010; // round
      10'b1100010001: out = 11'b10110011100;
      10'b1100010010: out = 11'b10110011111; // round
      10'b1100010011: out = 11'b10110100001; // round
      10'b1100010100: out = 11'b10110100011;
      10'b1100010101: out = 11'b10110100110; // round
      10'b1100010110: out = 11'b10110101000; // round
      10'b1100010111: out = 11'b10110101010;
      10'b1100011000: out = 11'b10110101101; // round
      10'b1100011001: out = 11'b10110101111;
      10'b1100011010: out = 11'b10110110001;
      10'b1100011011: out = 11'b10110110100; // round
      10'b1100011100: out = 11'b10110110110;
      10'b1100011101: out = 11'b10110111001; // round
      10'b1100011110: out = 11'b10110111011; // round
      10'b1100011111: out = 11'b10110111101;
      10'b1100100000: out = 11'b10111000000; // round
      10'b1100100001: out = 11'b10111000010;
      10'b1100100010: out = 11'b10111000101; // round
      10'b1100100011: out = 11'b10111000111; // round
      10'b1100100100: out = 11'b10111001001;
      10'b1100100101: out = 11'b10111001100; // round
      10'b1100100110: out = 11'b10111001110;
      10'b1100100111: out = 11'b10111010000;
      10'b1100101000: out = 11'b10111010011; // round
      10'b1100101001: out = 11'b10111010101;
      10'b1100101010: out = 11'b10111011000; // round
      10'b1100101011: out = 11'b10111011010;
      10'b1100101100: out = 11'b10111011100;
      10'b1100101101: out = 11'b10111011111; // round
      10'b1100101110: out = 11'b10111100001;
      10'b1100101111: out = 11'b10111100100; // round
      10'b1100110000: out = 11'b10111100110;
      10'b1100110001: out = 11'b10111101000;
      10'b1100110010: out = 11'b10111101011; // round
      10'b1100110011: out = 11'b10111101101;
      10'b1100110100: out = 11'b10111110000; // round
      10'b1100110101: out = 11'b10111110010;
      10'b1100110110: out = 11'b10111110101; // round
      10'b1100110111: out = 11'b10111110111; // round
      10'b1100111000: out = 11'b10111111001;
      10'b1100111001: out = 11'b10111111100; // round
      10'b1100111010: out = 11'b10111111110;
      10'b1100111011: out = 11'b11000000001; // round
      10'b1100111100: out = 11'b11000000011;
      10'b1100111101: out = 11'b11000000110; // round
      10'b1100111110: out = 11'b11000001000; // round
      10'b1100111111: out = 11'b11000001010;
      10'b1101000000: out = 11'b11000001101; // round
      10'b1101000001: out = 11'b11000001111;
      10'b1101000010: out = 11'b11000010010; // round
      10'b1101000011: out = 11'b11000010100;
      10'b1101000100: out = 11'b11000010111; // round
      10'b1101000101: out = 11'b11000011001; // round
      10'b1101000110: out = 11'b11000011011;
      10'b1101000111: out = 11'b11000011110; // round
      10'b1101001000: out = 11'b11000100000;
      10'b1101001001: out = 11'b11000100011; // round
      10'b1101001010: out = 11'b11000100101;
      10'b1101001011: out = 11'b11000101000; // round
      10'b1101001100: out = 11'b11000101010;
      10'b1101001101: out = 11'b11000101101; // round
      10'b1101001110: out = 11'b11000101111;
      10'b1101001111: out = 11'b11000110010; // round
      10'b1101010000: out = 11'b11000110100; // round
      10'b1101010001: out = 11'b11000110110;
      10'b1101010010: out = 11'b11000111001; // round
      10'b1101010011: out = 11'b11000111011;
      10'b1101010100: out = 11'b11000111110; // round
      10'b1101010101: out = 11'b11001000000;
      10'b1101010110: out = 11'b11001000011; // round
      10'b1101010111: out = 11'b11001000101;
      10'b1101011000: out = 11'b11001001000; // round
      10'b1101011001: out = 11'b11001001010;
      10'b1101011010: out = 11'b11001001101; // round
      10'b1101011011: out = 11'b11001001111;
      10'b1101011100: out = 11'b11001010010; // round
      10'b1101011101: out = 11'b11001010100;
      10'b1101011110: out = 11'b11001010111; // round
      10'b1101011111: out = 11'b11001011001;
      10'b1101100000: out = 11'b11001011100; // round
      10'b1101100001: out = 11'b11001011110;
      10'b1101100010: out = 11'b11001100001; // round
      10'b1101100011: out = 11'b11001100011;
      10'b1101100100: out = 11'b11001100110; // round
      10'b1101100101: out = 11'b11001101000;
      10'b1101100110: out = 11'b11001101011; // round
      10'b1101100111: out = 11'b11001101101;
      10'b1101101000: out = 11'b11001110000; // round
      10'b1101101001: out = 11'b11001110010;
      10'b1101101010: out = 11'b11001110101; // round
      10'b1101101011: out = 11'b11001110111;
      10'b1101101100: out = 11'b11001111010; // round
      10'b1101101101: out = 11'b11001111100;
      10'b1101101110: out = 11'b11001111111; // round
      10'b1101101111: out = 11'b11010000001;
      10'b1101110000: out = 11'b11010000100; // round
      10'b1101110001: out = 11'b11010000110;
      10'b1101110010: out = 11'b11010001001; // round
      10'b1101110011: out = 11'b11010001011;
      10'b1101110100: out = 11'b11010001110; // round
      10'b1101110101: out = 11'b11010010000;
      10'b1101110110: out = 11'b11010010011; // round
      10'b1101110111: out = 11'b11010010101;
      10'b1101111000: out = 11'b11010011000; // round
      10'b1101111001: out = 11'b11010011010;
      10'b1101111010: out = 11'b11010011101; // round
      10'b1101111011: out = 11'b11010011111;
      10'b1101111100: out = 11'b11010100010; // round
      10'b1101111101: out = 11'b11010100100;
      10'b1101111110: out = 11'b11010100111; // round
      10'b1101111111: out = 11'b11010101010; // round
      10'b1110000000: out = 11'b11010101100;
      10'b1110000001: out = 11'b11010101111; // round
      10'b1110000010: out = 11'b11010110001;
      10'b1110000011: out = 11'b11010110100; // round
      10'b1110000100: out = 11'b11010110110;
      10'b1110000101: out = 11'b11010111001; // round
      10'b1110000110: out = 11'b11010111011;
      10'b1110000111: out = 11'b11010111110; // round
      10'b1110001000: out = 11'b11011000000;
      10'b1110001001: out = 11'b11011000011;
      10'b1110001010: out = 11'b11011000110; // round
      10'b1110001011: out = 11'b11011001000;
      10'b1110001100: out = 11'b11011001011; // round
      10'b1110001101: out = 11'b11011001101;
      10'b1110001110: out = 11'b11011010000; // round
      10'b1110001111: out = 11'b11011010010;
      10'b1110010000: out = 11'b11011010101; // round
      10'b1110010001: out = 11'b11011011000; // round
      10'b1110010010: out = 11'b11011011010;
      10'b1110010011: out = 11'b11011011101; // round
      10'b1110010100: out = 11'b11011011111;
      10'b1110010101: out = 11'b11011100010; // round
      10'b1110010110: out = 11'b11011100100;
      10'b1110010111: out = 11'b11011100111; // round
      10'b1110011000: out = 11'b11011101010; // round
      10'b1110011001: out = 11'b11011101100;
      10'b1110011010: out = 11'b11011101111; // round
      10'b1110011011: out = 11'b11011110001;
      10'b1110011100: out = 11'b11011110100; // round
      10'b1110011101: out = 11'b11011110111; // round
      10'b1110011110: out = 11'b11011111001;
      10'b1110011111: out = 11'b11011111100; // round
      10'b1110100000: out = 11'b11011111110;
      10'b1110100001: out = 11'b11100000001; // round
      10'b1110100010: out = 11'b11100000011;
      10'b1110100011: out = 11'b11100000110;
      10'b1110100100: out = 11'b11100001001; // round
      10'b1110100101: out = 11'b11100001011;
      10'b1110100110: out = 11'b11100001110; // round
      10'b1110100111: out = 11'b11100010001; // round
      10'b1110101000: out = 11'b11100010011;
      10'b1110101001: out = 11'b11100010110; // round
      10'b1110101010: out = 11'b11100011000;
      10'b1110101011: out = 11'b11100011011; // round
      10'b1110101100: out = 11'b11100011110; // round
      10'b1110101101: out = 11'b11100100000;
      10'b1110101110: out = 11'b11100100011; // round
      10'b1110101111: out = 11'b11100100101;
      10'b1110110000: out = 11'b11100101000;
      10'b1110110001: out = 11'b11100101011; // round
      10'b1110110010: out = 11'b11100101101;
      10'b1110110011: out = 11'b11100110000; // round
      10'b1110110100: out = 11'b11100110011; // round
      10'b1110110101: out = 11'b11100110101;
      10'b1110110110: out = 11'b11100111000; // round
      10'b1110110111: out = 11'b11100111011; // round
      10'b1110111000: out = 11'b11100111101;
      10'b1110111001: out = 11'b11101000000; // round
      10'b1110111010: out = 11'b11101000010;
      10'b1110111011: out = 11'b11101000101;
      10'b1110111100: out = 11'b11101001000; // round
      10'b1110111101: out = 11'b11101001010;
      10'b1110111110: out = 11'b11101001101;
      10'b1110111111: out = 11'b11101010000; // round
      10'b1111000000: out = 11'b11101010010;
      10'b1111000001: out = 11'b11101010101; // round
      10'b1111000010: out = 11'b11101011000; // round
      10'b1111000011: out = 11'b11101011010;
      10'b1111000100: out = 11'b11101011101; // round
      10'b1111000101: out = 11'b11101100000; // round
      10'b1111000110: out = 11'b11101100010;
      10'b1111000111: out = 11'b11101100101; // round
      10'b1111001000: out = 11'b11101101000; // round
      10'b1111001001: out = 11'b11101101010;
      10'b1111001010: out = 11'b11101101101; // round
      10'b1111001011: out = 11'b11101110000; // round
      10'b1111001100: out = 11'b11101110010;
      10'b1111001101: out = 11'b11101110101;
      10'b1111001110: out = 11'b11101111000; // round
      10'b1111001111: out = 11'b11101111010;
      10'b1111010000: out = 11'b11101111101;
      10'b1111010001: out = 11'b11110000000; // round
      10'b1111010010: out = 11'b11110000010;
      10'b1111010011: out = 11'b11110000101;
      10'b1111010100: out = 11'b11110001000; // round
      10'b1111010101: out = 11'b11110001010;
      10'b1111010110: out = 11'b11110001101;
      10'b1111010111: out = 11'b11110010000; // round
      10'b1111011000: out = 11'b11110010011; // round
      10'b1111011001: out = 11'b11110010101;
      10'b1111011010: out = 11'b11110011000; // round
      10'b1111011011: out = 11'b11110011011; // round
      10'b1111011100: out = 11'b11110011101;
      10'b1111011101: out = 11'b11110100000;
      10'b1111011110: out = 11'b11110100011; // round
      10'b1111011111: out = 11'b11110100110; // round
      10'b1111100000: out = 11'b11110101000;
      10'b1111100001: out = 11'b11110101011; // round
      10'b1111100010: out = 11'b11110101110; // round
      10'b1111100011: out = 11'b11110110000;
      10'b1111100100: out = 11'b11110110011;
      10'b1111100101: out = 11'b11110110110; // round
      10'b1111100110: out = 11'b11110111001; // round
      10'b1111100111: out = 11'b11110111011;
      10'b1111101000: out = 11'b11110111110; // round
      10'b1111101001: out = 11'b11111000001; // round
      10'b1111101010: out = 11'b11111000011;
      10'b1111101011: out = 11'b11111000110;
      10'b1111101100: out = 11'b11111001001; // round
      10'b1111101101: out = 11'b11111001100; // round
      10'b1111101110: out = 11'b11111001110;
      10'b1111101111: out = 11'b11111010001;
      10'b1111110000: out = 11'b11111010100; // round
      10'b1111110001: out = 11'b11111010111; // round
      10'b1111110010: out = 11'b11111011001;
      10'b1111110011: out = 11'b11111011100;
      10'b1111110100: out = 11'b11111011111; // round
      10'b1111110101: out = 11'b11111100010; // round
      10'b1111110110: out = 11'b11111100100;
      10'b1111110111: out = 11'b11111100111;
      10'b1111111000: out = 11'b11111101010; // round
      10'b1111111001: out = 11'b11111101101; // round
      10'b1111111010: out = 11'b11111101111;
      10'b1111111011: out = 11'b11111110010;
      10'b1111111100: out = 11'b11111110101; // round
      10'b1111111101: out = 11'b11111111000; // round
      10'b1111111110: out = 11'b11111111010;
      10'b1111111111: out = 11'b11111111101;
      default: out = 11'bxxxxxxxxxxx;
    endcase
  end
endmodule
