// Copyright (c) Facebook, Inc. and its affiliates. All Rights Reserved.
// All rights reserved.
//
// This source code is licensed under the license found in the
// LICENSE file in the root directory of this source tree.


//
// (8, 1)-log
//

// how large the CPU wrapper size is
parameter CONFIG_LOG_WRAP_BITS = 8;
parameter CONFIG_LOG_WIDTH = 8;
parameter CONFIG_LOG_LS = 1;
parameter CONFIG_LOG_TO_LINEAR_BITS = 5;
parameter CONFIG_LINEAR_TO_LOG_BITS = 5;

parameter CONFIG_LOG_ACC_WRAP_BITS = 64;
parameter CONFIG_LOG_ACC_BITS = 41;
